library verilog;
use verilog.vl_types.all;
entity tb_Pipeline is
end tb_Pipeline;
