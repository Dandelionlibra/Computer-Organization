// 設定時間尺度
`timescale 1ns/1ns
// 定義 module ID_EX 可連接的 ports
module ID_EX( clk, reset, next_PC_ID, );
// 定義哪些 ports 為 input，哪些為 output
input clk;
input reset;



endmodule