// 設定時間尺度
`timescale 1ns/1ns
// 定義 module EX_MEM 可連接的 ports
module EX_MEM( clk, reset, , MenRW_EX, MenRW_MEM, Branch_EX, Branch_MEM );
// 定義哪些 ports 為 input，哪些為 output
input clk;
input reset;



endmodule